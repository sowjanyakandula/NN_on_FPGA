`timescale 1ns / 1ps

module weight_read_testbench();
   reg clk,rst;
   wire [7:0] dout;
   wire [7:0] dummy;
   wire [11:0] wout;
   integer f,i;

  
 
   
 
   
endmodule