`timescale 1ns / 1ps

module pro_multi(
    input [31:0] A,
    input [31:0] B,
    output [31:0] Res,
    input clk
    );
    
endmodule
