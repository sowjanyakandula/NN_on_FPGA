`timescale 1ns / 1ps

module test_bench_final_code();
    reg clk,rst;
   wire [7:0] dout;
   integer f,i;

  

endmodule
